** Profile: "SCHEMATIC1-CA1-Q2-D-Current_Source-Simulate"  [ E:\UT Programming\Electrical-Circuits-Fall-2024\CA1\Q2\D\Current Source\ca1-q2-d-current_source-SCHEMATIC1-CA1-Q2-D-Current_Source-Simulate.sim ] 

** Creating circuit file "ca1-q2-d-current_source-SCHEMATIC1-CA1-Q2-D-Current_Source-Simulate.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN I_I1 0 10 0.5 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\ca1-q2-d-current_source-SCHEMATIC1.net" 


.END
