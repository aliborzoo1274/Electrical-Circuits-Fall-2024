** Profile: "SCHEMATIC1-Q1-Simulate"  [ E:\UT Programming\Electrical-Circuits-Fall-2024\CA1\ca1-q1-schematic1-q1-simulate.sim ] 

** Creating circuit file "ca1-q1-schematic1-q1-simulate.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\ca1-q1-SCHEMATIC1.net" 


.END
