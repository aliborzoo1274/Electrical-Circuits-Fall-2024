** Profile: "SCHEMATIC1-CA1-Q3-B-Simulate"  [ E:\UT Programming\Electrical-Circuits-Fall-2024\CA1\Q3\B\ca1-q3-b-schematic1-ca1-q3-b-simulate.sim ] 

** Creating circuit file "ca1-q3-b-schematic1-ca1-q3-b-simulate.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\ca1-q3-b-SCHEMATIC1.net" 


.END
