** Profile: "SCHEMATIC1-CA1-Q3-C-Simulate"  [ E:\UT Programming\Electrical-Circuits-Fall-2024\CA1\Q3\C\ca1-q3-c-SCHEMATIC1-CA1-Q3-C-Simulate.sim ] 

** Creating circuit file "ca1-q3-c-SCHEMATIC1-CA1-Q3-C-Simulate.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN PARAM RLval 0.5 50 0.5 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\ca1-q3-c-SCHEMATIC1.net" 


.END
