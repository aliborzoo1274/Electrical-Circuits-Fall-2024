** Profile: "SCHEMATIC1-CA1-Q2-A-Simulate"  [ E:\UT PROGRAMMING\ELECTRICAL-CIRCUITS-FALL-2024\CA1\Q2\A\ca1-q2-a-SCHEMATIC1-CA1-Q2-A-Simulate.sim ] 

** Creating circuit file "ca1-q2-a-SCHEMATIC1-CA1-Q2-A-Simulate.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\ca1-q2-a-SCHEMATIC1.net" 


.END
