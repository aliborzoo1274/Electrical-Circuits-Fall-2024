** Profile: "SCHEMATIC1-CA1-Q3-D-Simulate"  [ E:\UT Programming\Electrical-Circuits-Fall-2024\CA1\Q3\D\ca1-q3-d-SCHEMATIC1-CA1-Q3-D-Simulate.sim ] 

** Creating circuit file "ca1-q3-d-SCHEMATIC1-CA1-Q3-D-Simulate.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 10ms 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\ca1-q3-d-SCHEMATIC1.net" 


.END
