** Profile: "SCHEMATIC1-CA1-Q2-D-Voltage_Source"  [ E:\UT Programming\Electrical-Circuits-Fall-2024\CA1\Q2\D\Voltage Source\ca1-q2-d-voltage_source-SCHEMATIC1-CA1-Q2-D-Voltage_Source.sim ] 

** Creating circuit file "ca1-q2-d-voltage_source-SCHEMATIC1-CA1-Q2-D-Voltage_Source.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN V_V1 0 10 0.5 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\ca1-q2-d-voltage_source-SCHEMATIC1.net" 


.END
